`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06.04.2025 15:38:08
// Design Name: 
// Module Name: 
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
//Function 1 is Normalizing
//Function 2 is Rounding
/*
Normalizing unit:
inputs: 112 bit long mantissa
11 bit long exponent
1 bit sign
2 bit opcode
*/
module norm_rnd (clk, fract_in, exp_in, sign, opcode, remainder, r_mode,
                fract_out, exp_out, dn_out, ine_out, overflow_out, infinite_out);
    input clk;
    input [105:0] fract_in;
    input [10:0] exp_in;
    input sign; //Rounding only
    input [1:0] opcode; //Rounding only
    input [52:0] remainder; //Rounding only
    input [1:0] r_mode; //Rounding only
    
    output reg [52:0] fract_out;
    output reg [10:0] exp_out;
    output reg dn_out;
    output reg ine_out;
    output reg overflow_out;
    output reg infinite_out;
                

    //Local Wires & Registers
    reg [6:0] fract_1dz;    /*reg needed to hold the value constantly - register should not be clocked as it is fed by
                            combi circuit - up to 111 leading zeros may be present, thus
                            a 7 bit register is needed*/
    wire shift_dir;         //Direction of shift
    wire exp_max;           //Exponent is max
    wire [6:0] shift_val;   //Magnitude of shift
    wire ldz_less_exp;      //Exponent is larger than no of left shifts required
    wire [6:0] fract_1dz_nil;
    wire [10:0] exp_in_nil;
    wire out_dn;            //indicates that the outputwillbe denormalized
    wire out_overflow;      //indicates that output overflow occured- exponent& mantissa cannot store result
    wire [105:0] fract_sh_R, fract_sh_L;
    wire [10:0] exp_sh_R, exp_sh_L;
    wire [105:0] fract_shifted;
    wire [10:0] exp_shifted;
    
    wire [52:0] fract_down, fract_up_temp,fract_up; //wireto store rounded down&up fractions
    wire cout;                                      //wire to store carry out from fractjip
    wire [10:0] exp_up;                             //wire to store exponent for fractjip - 
                                                    //needed becoz fractjip may have carry-out
    wire fract_trunc;                                //indicates that some value have been truncated
    wire rem_not_zero;                              //indicates that the division has a non-zero remainder- 
                                                    //used to signal inexact
                                                    
    reg [52:0] fract_round;
    reg [10:0] exp_round;
    wire [52:0] fract_near_temp, fract_round_nearest, fract_round_zero; //stores result for every rounding mode
    reg [52:0] fract_round_up, fract_round_down; //stores result for every rounding mode
    wire [10:0] exp_near_temp, exp_round_nearest, exp_round_zero;
    reg [10:0] exp_round_up, exp_round_down;
    wire last_bit, trunc, r_near_sel, fract_up_overflow;
    wire [1:0] r_up_sel, r_down_sel;
    
    always @ (fract_in)
        casex (fract_in) // synopsys full_case parallel_case
            106'b1?????????????????????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 0;
            106'b01????????????????????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 1;
            106'b001???????????????????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 2;
            106'b0001??????????????????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 3;
            106'b00001?????????????????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 4;
            106'b000001????????????????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 5;
            106'b0000001???????????????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 6;
            106'b00000001??????????????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 7;
            106'b000000001?????????????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 8;
            106'b0000000001????????????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 9;
            106'b00000000001???????????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 10;
            106'b000000000001??????????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 11;
            106'b0000000000001?????????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 12;
            106'b00000000000001????????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 13;
            106'b000000000000001???????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 14;
            106'b0000000000000001??????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 15;
            106'b00000000000000001?????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 16;
            106'b000000000000000001????????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 17;
            106'b0000000000000000001???????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 18;
            106'b00000000000000000001??????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 19;
            106'b000000000000000000001?????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 20;
            106'b0000000000000000000001????????????????????????????????????????????????????????????????????????????????????: fract_1dz = 21;
            106'b00000000000000000000001???????????????????????????????????????????????????????????????????????????????????: fract_1dz = 22;
            106'b000000000000000000000001??????????????????????????????????????????????????????????????????????????????????: fract_1dz = 23;
            106'b0000000000000000000000001?????????????????????????????????????????????????????????????????????????????????: fract_1dz = 24;
            106'b00000000000000000000000001????????????????????????????????????????????????????????????????????????????????: fract_1dz = 25;
            106'b000000000000000000000000001???????????????????????????????????????????????????????????????????????????????: fract_1dz = 26;
            106'b0000000000000000000000000001??????????????????????????????????????????????????????????????????????????????: fract_1dz = 27;
            106'b00000000000000000000000000001?????????????????????????????????????????????????????????????????????????????: fract_1dz = 28;
            106'b000000000000000000000000000001????????????????????????????????????????????????????????????????????????????: fract_1dz = 29;
            106'b0000000000000000000000000000001???????????????????????????????????????????????????????????????????????????: fract_1dz = 30;
            106'b00000000000000000000000000000001??????????????????????????????????????????????????????????????????????????: fract_1dz = 31;
            106'b000000000000000000000000000000001?????????????????????????????????????????????????????????????????????????: fract_1dz = 32;
            106'b0000000000000000000000000000000001????????????????????????????????????????????????????????????????????????: fract_1dz = 33;
            106'b00000000000000000000000000000000001???????????????????????????????????????????????????????????????????????: fract_1dz = 34;
            106'b000000000000000000000000000000000001??????????????????????????????????????????????????????????????????????: fract_1dz = 35;
            106'b0000000000000000000000000000000000001?????????????????????????????????????????????????????????????????????: fract_1dz = 36;
            106'b00000000000000000000000000000000000001????????????????????????????????????????????????????????????????????: fract_1dz = 37;
            106'b000000000000000000000000000000000000001???????????????????????????????????????????????????????????????????: fract_1dz = 38;
            106'b0000000000000000000000000000000000000001??????????????????????????????????????????????????????????????????: fract_1dz = 39;
            106'b00000000000000000000000000000000000000001?????????????????????????????????????????????????????????????????: fract_1dz = 40;
            106'b000000000000000000000000000000000000000001????????????????????????????????????????????????????????????????: fract_1dz = 41;
            106'b0000000000000000000000000000000000000000001???????????????????????????????????????????????????????????????: fract_1dz = 42;
            106'b00000000000000000000000000000000000000000001??????????????????????????????????????????????????????????????: fract_1dz = 43;
            106'b000000000000000000000000000000000000000000001?????????????????????????????????????????????????????????????: fract_1dz = 44;
            106'b0000000000000000000000000000000000000000000001????????????????????????????????????????????????????????????: fract_1dz = 45;
            106'b00000000000000000000000000000000000000000000001???????????????????????????????????????????????????????????: fract_1dz = 46;
            106'b000000000000000000000000000000000000000000000001??????????????????????????????????????????????????????????: fract_1dz = 47;
            106'b0000000000000000000000000000000000000000000000001?????????????????????????????????????????????????????????: fract_1dz = 48;
            106'b00000000000000000000000000000000000000000000000001????????????????????????????????????????????????????????: fract_1dz = 49;
            106'b000000000000000000000000000000000000000000000000001???????????????????????????????????????????????????????: fract_1dz = 50;
            106'b0000000000000000000000000000000000000000000000000001??????????????????????????????????????????????????????: fract_1dz = 51;
            106'b00000000000000000000000000000000000000000000000000001?????????????????????????????????????????????????????: fract_1dz = 52;
            106'b000000000000000000000000000000000000000000000000000001????????????????????????????????????????????????????: fract_1dz = 53;
            106'b0000000000000000000000000000000000000000000000000000001???????????????????????????????????????????????????: fract_1dz = 54;
            106'b00000000000000000000000000000000000000000000000000000001??????????????????????????????????????????????????: fract_1dz = 55;
            106'b000000000000000000000000000000000000000000000000000000001?????????????????????????????????????????????????: fract_1dz = 56;
            106'b0000000000000000000000000000000000000000000000000000000001????????????????????????????????????????????????: fract_1dz = 57;
            106'b00000000000000000000000000000000000000000000000000000000001???????????????????????????????????????????????: fract_1dz = 58;
            106'b000000000000000000000000000000000000000000000000000000000001??????????????????????????????????????????????: fract_1dz = 59;
            106'b0000000000000000000000000000000000000000000000000000000000001?????????????????????????????????????????????: fract_1dz = 60;
            106'b00000000000000000000000000000000000000000000000000000000000001????????????????????????????????????????????: fract_1dz = 61;
            106'b000000000000000000000000000000000000000000000000000000000000001???????????????????????????????????????????: fract_1dz = 62;
            106'b0000000000000000000000000000000000000000000000000000000000000001??????????????????????????????????????????: fract_1dz = 63;
            106'b00000000000000000000000000000000000000000000000000000000000000001?????????????????????????????????????????: fract_1dz = 64;
            106'b000000000000000000000000000000000000000000000000000000000000000001????????????????????????????????????????: fract_1dz = 65;
            106'b0000000000000000000000000000000000000000000000000000000000000000001???????????????????????????????????????: fract_1dz = 66;
            106'b00000000000000000000000000000000000000000000000000000000000000000001??????????????????????????????????????: fract_1dz = 67;
            106'b000000000000000000000000000000000000000000000000000000000000000000001?????????????????????????????????????: fract_1dz = 68;
            106'b0000000000000000000000000000000000000000000000000000000000000000000001????????????????????????????????????: fract_1dz = 69;
            106'b00000000000000000000000000000000000000000000000000000000000000000000001???????????????????????????????????: fract_1dz = 70;
            106'b000000000000000000000000000000000000000000000000000000000000000000000001??????????????????????????????????: fract_1dz = 71;
            106'b0000000000000000000000000000000000000000000000000000000000000000000000001?????????????????????????????????: fract_1dz = 72;
            106'b00000000000000000000000000000000000000000000000000000000000000000000000001????????????????????????????????: fract_1dz = 73;
            106'b000000000000000000000000000000000000000000000000000000000000000000000000001???????????????????????????????: fract_1dz = 74;
            106'b0000000000000000000000000000000000000000000000000000000000000000000000000001??????????????????????????????: fract_1dz = 75;
            106'b00000000000000000000000000000000000000000000000000000000000000000000000000001?????????????????????????????: fract_1dz = 76;
            106'b000000000000000000000000000000000000000000000000000000000000000000000000000001????????????????????????????: fract_1dz = 77;
            106'b0000000000000000000000000000000000000000000000000000000000000000000000000000001???????????????????????????: fract_1dz = 78;
            106'b00000000000000000000000000000000000000000000000000000000000000000000000000000001??????????????????????????: fract_1dz = 79;
            106'b000000000000000000000000000000000000000000000000000000000000000000000000000000001?????????????????????????: fract_1dz = 80;
            106'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001????????????????????????: fract_1dz = 81;
            106'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001???????????????????????: fract_1dz = 82;
            106'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001??????????????????????: fract_1dz = 83;
            106'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001?????????????????????: fract_1dz = 84;
            106'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001????????????????????: fract_1dz = 85;
            106'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001???????????????????: fract_1dz = 86;
            106'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001??????????????????: fract_1dz = 87;
            106'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001?????????????????: fract_1dz = 88;
            106'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001????????????????: fract_1dz = 89;
            106'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001???????????????: fract_1dz = 90;
            106'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001??????????????: fract_1dz = 91;
            106'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001?????????????: fract_1dz = 92;
            106'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001????????????: fract_1dz = 93;
            106'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001???????????: fract_1dz = 94;
            106'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001??????????: fract_1dz = 95;
            106'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001?????????: fract_1dz = 96;
            106'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001????????: fract_1dz = 97;
            106'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001???????: fract_1dz = 98;
            106'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001??????: fract_1dz = 99;
            106'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001?????: fract_1dz = 100;
            106'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001????: fract_1dz = 101;
            106'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001???: fract_1dz = 102;
            106'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001??: fract_1dz = 103;
            106'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001?: fract_1dz = 104;
            106'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: fract_1dz = 105;
        endcase
        
    assign shift_dir= -(|fract_1dz); //shift_dir - 0 meansleft,shiftjiir = 1meansright
    assign exp_max = &exp_in[10:1];
    assign ldz_less_exp = (fract_1dz <= exp_in[6:0]) ? 1'b1 : |exp_in[10:7];
    assign fract_1dz_nil = fract_1dz -1;
    assign exp_in_nil = exp_in - 1;
    assign shift_val = ldz_less_exp ? fract_1dz_nil : exp_in_nil;
    
    assign fract_sh_R = fract_in >> 1'b1;
    assign exp_sh_R = exp_in + 1;
    assign fract_sh_L = fract_in << shift_val;
    assign exp_sh_L = exp_in - shift_val;
    
    assign fract_shifted = (fract_1dz == 1)? fract_in : (shift_dir) ? fract_sh_R: fract_sh_L;
    assign exp_shifted = (fract_1dz == 1) ? (exp_in): ((shift_dir) ? exp_sh_R : exp_sh_L );
    
    assign out_dn = !ldz_less_exp;
    assign out_overflow = (exp_max & shift_dir);
    
    //rounded
    assign fract_down = fract_shifted[104:52];
    assign {cout, fract_up_temp} = fract_down + {53'b0, 1'b1};
    
    assign fract_up = (cout)? {cout, fract_up_temp} >> 1 : fract_up_temp;
    assign exp_up = exp_shifted + {10'b0,cout};
    assign fract_up_overflow = cout & (&exp_shifted[10:1]);
    
    assign lastbit = fract_shifted[51];
    
    assign trunc = |fract_shifted[50:0];
    
    assign r_near_sel= last_bit & (trunc | fract_down[0]); 
    
    assign fract_near_temp = (r_near_sel) ? fract_up : fract_down;
    
    assign exp_near_temp = (r_near_sel) ? exp_up : exp_shifted;
    
    assign fract_round_nearest = (out_overflow | (r_near_sel & fract_up_overflow)) ? 53'b0 : fract_near_temp;
    
    assign exp_round_nearest = (out_overflow | (r_near_sel & fract_up_overflow)) ? 11'h7FF : exp_near_temp;
    
    //Round to zero calculation
    assign fract_round_zero = (out_overflow) ? 53'h1FFFFFFFFFFFFF : fract_down;
    assign exp_round_ero = (out_overflow) ? 11'h7FE: exp_shifted;

    //Round up calculation
    assign r_up_sel[0] = sign;
    assign r_up_sel[1] = out_overflow | (-sign &fract_up_overflow);
    
    always @(r_up_sel or fract_up or fract_down)
        case (r_up_sel)
            2'b00 : fract_round_up = fract_up;
            2'b01 : fract_round_up = fract_up;
            2'b10 : fract_round_up = 53'b0;
            2'b11 : fract_round_up = 53'h1FFFFFFFFFFFFF;
        endcase
        
    always @(r_up_sel or exp_up or exp_shifted)
        case (r_up_sel) // synopsys full_caseparallelj;ase
            2'b00 : exp_round_up = exp_up;
            2'b01 : exp_round_up = exp_shifted;
            2'b10 : exp_round_up = 11'h7FF;
            2'b11 : exp_round_up = 11'h7FE;
        endcase
        
        assign r_down_sel[0] = -sign;
        assign r_down_sel[1] = out_overflow | (sign & fract_up_overflow);
        always @(r_down_sel or fract_up or fract_down)
            case (r_down_sel) // synopsys full_caseparallel_case
            2'b00 : fract_round_down = fract_up;
            2'b01 : fract_round_down = fract_down;
            2'b10 : fract_round_down = 53'b0;
            2'b11 : fract_round_down = 53'h1FFFFFFFFFFFFF;
        endcase
        
        always @(r_down_sel or exp_up or exp_shifted)
            case (r_down_sel) // synopsys full_case parallel_case
            2'b00 : exp_round_down = exp_up;
            2'b01 : exp_round_down = exp_shifted;
            2'b10 : exp_round_down = 11'h7FF;
            2'b11 : exp_round_down = 11'h7FE;
        endcase
    
    always @(r_mode or fract_round_nearest or fract_round_zero or fract_round_up or fract_round_down)
        case (r_mode)
            2'b00 : fract_round = fract_round_nearest;
            2'b01 : fract_round = fract_round_zero;
            2'b10 : fract_round = fract_round_up;
            2'b11 : fract_round = fract_round_down;
        endcase
    
    always @(r_mode or fract_round_nearest or fract_round_zero or fract_round_up or fract_round_down)
        case (r_mode)
            2'b00 : exp_round = exp_round_nearest;
            2'b01 : exp_round = exp_round_zero;
            2'b10 : exp_round = exp_round_up;
            2'b11 : exp_round = exp_round_down;
        endcase
        
    assign fract_trunc = last_bit | trunc;
    assign rem_not_zero = (&opcode) & (|remainder);
    
    always @(posedge clk)
        begin
            fract_out <= fract_round;
            exp_out <= exp_round;
            dn_out <= out_dn;
            ine_out <= fract_trunc | rem_not_zero;
            overflow_out <= out_overflow;
            infinite_out <= out_overflow &((|r_mode)|(r_mode[1] & ~(r_mode[0]^sign)));
        end
        
       
    
    
endmodule